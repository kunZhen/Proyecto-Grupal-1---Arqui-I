module Bilinea(
	input logic clk, reset
	
);

endmodule 