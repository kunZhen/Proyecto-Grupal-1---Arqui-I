module PISA(
	input logic clk, reset
	
);
	

endmodule 